import axi_helper::*;
module subordinate(	
	axi4_if.subordinate_mp bus,
	TB_if.subordinate tb
	);
	localparam DATA_W = axi4_if.DATA_W;				//pull in DATA_W
	localparam ADDR_W = axi4_if.ADDR_W;				//pull in ADDR_W
	byte unsigned memory [0:4095];				//cache is smaller than memory! CPU
	logic [DATA_W:0] data_W, data_R;			  	//data_W,addr_AW,addr_R, opcode
	logic [ADDR_W:0] addr_AW, addr_AR;				//hook input address for AW 
								
	logic [4:0] rx_flag,tx_flag;				//data flag register notifies if new data present on channel latch (if RX
	
	logic zero,bresp; 
	
	resp_t tx_bresp, tx_rresp;
	assign tx_bresp = OKAY;					//these are hanging ports for now
	assign tx_rresp = OKAY;
	assign zero  = 1'b0;
	
	/*============= AW CHANNEL =============*/
	RX_channel AW #(.WIDTH(ADDR_W))(				//Write DATA
		.ACLK(bus.ACLK),
		.ARESETn(bus.ARESETn),						
	 	.READY(bus.AWREADY),
		.VALID(bus.AWVALID),
		.xDATA(bus.AWDATA),
		
		.rx_data(tb.sub_rx_AW),				//DATA RECIEVED BY SUB	
	 	.rx_new_data(tb.new_data[4]),			//flag for new data recieved
		.rx_hold(tb.mem_flag[4]),				//1: SUB says HOLD the transfer for processing
	);
	/*============= W CHANNEL =============*/
	RX_channel W #(.WIDTH(DATA_W))(				//Write DATA	
		.ACLK(bus.ACLK),
		.ARESETn(bus.ARESETn),						
	 	.READY(bus.WREADY),
		.VALID(bus.WVALID),
		.xDATA(bus.WDATA),
		
		.rx_data(tb.sub_rx_W),						
	 	.rx_new_data(tb.new_data[3]),			
		.rx_hold(tb.mem_flag[3]),
	);
	/*============= B CHANNEL =============*/
	TX_channel B #(.WIDTH(2))(				//write confirmation channel B
		.ACLK(bus.ACLK),
		.ARESETn(bus.ARESETn),						
	 	.READY(bus.BREADY),
	 	.VALID(bus.BVALID),
	 	.xDATA(bus.BDATA),
	 	
	 	.tx_data(rb.sub_bresp),
	 	.tx_en(tb.tx_en[2]),
	 	.tx_hold()				
	);	
	/*============= AR CHANNEL =============*/
	RX_channel AR #(.WIDTH(ADDR_W))(				//READ address DATA
		.ACLK(bus.ACLK),
		.ARESETn(bus.ARESETn),						
	 	.READY(bus.ARREADY),
		.VALID(bus.ARVALID),
		.xDATA(bus.ARDATA),
		
		.rx_data(tb.sub_rx_AR),				
	 	.rx_new_data(tb.new_data[1]),			
		.rx_hold(tb.mem_flag[1]),
	);
	/*============= R CHANNEL =============*/
	TX_channel R #(.WIDTH(DATA_W))(				//Read channel 
		.ACLK(bus.ACLK),
		.ARESETn(bus.ARESETn),						
	 	.READY(bus.RREADY),
	 	.VALID(bus.RVALID),
	 	.xDATA(bus.RDATA),
	 	
	 	.tx_data(tb.sub_tx_R),				//outgoing data from SUB
	 	.tx_en(tb.tx_en[0]),				//SUB enables the transfer
	 	.tx_hold()					//~READY from the master use this or (~bus.RREADY)
	);
	
	//reset is handled in RX/TX modules where states are set to idle Valid = 0/ready =1
	

endmodule

/* 
	always_comb begin 
		bresp = 2'b00;
		AWW_latched = data_flag[4] & data_flag[3];
		if (data_flag[1]) begin
			data_R = memory [addr_AR];			//asynchronous read
		end
	end
	always_ff @ (posedge ACLK) begin 
		if (ARESETn)
		else

	end
*/
/*
	Mem_Manager_Write R_service #(
		.LEN_ADDR(12),
		.LEN_DATA(DATA_W) 
		)(							//master has 11 addr and slave has 10, cs of which slave is the 11th address
		.*,							//aCLK,ARESETn,
		.ADDR(addr_AW[11:0]),					//take the bottom 32 bit→ SET/INDEX we'll just overwirte data in cache
		.DATA(data_R),
		.WE(.data_flag[0]), 					//write enable
		.memory(memory),					//*** passes whole memory maybe better to pass by refference?
		.MEM_BUSY(mem_flag[0])
	);
*/
